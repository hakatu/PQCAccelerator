//////////////////////////////////////////////////////////////////////////////////
//
//
// Filename        : compute_unit.sv
// Description     : Compute unit main branches 4 FIFO 2 input Compute Core
//
//////////////////////////////////////////////////////////////////////////////////

module compute_unit (
    clk,
    rst,

    //usage interface 
    idat1,
    idat2,
    idatwr,
    inrdy, //rdy take input


    odat1,
    odat2,
    odatrd,
    outrdy, //rdy take output
    //////
)


////////////generate 4 FF circle


endmodule